class env_config;
 virtual tinyalu_bfm bfm;

 function new(virtual tinyalu_bfm bfm);
    this.bfm = bfm;
 endfunction : new
 
endclass : env_config

