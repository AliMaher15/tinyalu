interface tinyalu_bfm;

  // import pakage
  import tinyalu_pkg::*;
  
  // variables declaration
  byte         unsigned        A;
  byte         unsigned        B;
  bit          clk;
  bit          reset_n;
  wire [2:0]   op;
  bit          start;
  wire         done;
  wire [15:0]  result;
  operation_t  op_set; 

  // monitors handles
  command_monitor command_monitor_h;
  result_monitor  result_monitor_h;

  assign op = op_set;

  task reset_alu();
    reset_n = 1'b0;  // activate
    @(negedge clk);
    @(negedge clk);
    reset_n = 1'b1; // deactivate
    start = 1'b0;
  endtask : reset_alu

  task send_op(input byte iA, input byte iB, input operation_t iop, output shortint alu_result);
    if (iop == rst_op) begin // rst op
      @(posedge clk);
      reset_n = 1'b0; // activate
      start = 1'b0;
      @(posedge clk);
      #1; // just to be sure
      reset_n = 1'b1; // deactivate
    end else begin // other 
      @(negedge clk);
      op_set = iop;
      A = iA;
      B = iB;
      start = 1'b1;
      if (iop == no_op) begin // no op
        @(posedge clk);
        #1;
        start = 1'b0;
      end else begin // add~mul
        do
          @(negedge clk); // loop to wait for operation to finish
        while (done == 0);
        alu_result = result;
        start = 1'b0; // done
      end
    end // else: !if(iop == rst_op)
  endtask : send_op

  function operation_t op2enum();
    case (op)
      3'b000 : return no_op;
      3'b001 : return add_op;
      3'b010 : return and_op;
      3'b011 : return xor_op;
      3'b100 : return mul_op;
      default : $fatal("Illegal operation on op bus");
    endcase
  endfunction : op2enum
  
  always @(posedge clk) begin : op_monitor
   static bit in_command = 0;
   if (start) begin : start_high
      if(!in_command) begin : new_command
        command_monitor_h.write_to_monitor(A, B, op2enum()); //send input to input monitor
        in_command = (op2enum() != no_op); // if no_op then no new command "0"
      end : new_command
    end : start_high
    else // start low
      in_command = 0;
  end : op_monitor

  // I am not sure about this always (its meaning)
  always @(negedge reset_n) begin : rst_monitor
    if (command_monitor_h != null) //guard against VCS time 0 negedge
       command_monitor_h.write_to_monitor($random,0,rst_op);
  end : rst_monitor  

  initial begin : result_monitor_thread
     forever begin : result_monitor_block
        @(posedge clk) ;
        if (done) 
          result_monitor_h.write_to_monitor(result); // send o/p when done
     end : result_monitor_block
  end : result_monitor_thread

  initial begin // clock generation
    clk = 0;
    fork
      forever begin
        #10
        clk = ~clk;
      end
    join_none
  end

endinterface : tinyalu_bfm